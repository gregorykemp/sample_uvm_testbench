// ----------------------------------------
// Wrapper object for test configuration.

class my_config extends uvm_object;

   int num_tx;

endclass : my_config