// ------------------------------------------------------------------------------
// Define UVM testbench package.

// Import UVM packages.
import uvm_pkg::*;

package vscale_mul_div_pkg;

   // Include UVM macros 
   `include "uvm_macros.svh"

   // Include testbench components and objects
   

endpackage : vscale_mul_div_pkg